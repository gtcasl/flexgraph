module fp_mult (
		input  wire [31:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire [31:0] b,      //      b.b
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [31:0] q       //      q.q
	);
endmodule

